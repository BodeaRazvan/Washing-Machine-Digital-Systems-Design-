library IEEE;
use IEEE.STD_LOGIC_1164.all; 
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ROM_WASH is	 
	port(
	I:in std_logic_vector (18 downto 0);
	Z:out std_logic_vector (35 downto 0)
	);
end ROM_WASH;



architecture ROM_WASH of ROM_WASH is  
type mem is array(0 to 818) of std_logic_vector (35 downto 0);
constant values :mem:=(	
x"000000000",
x"045304000",
x"145304000",
x"222302000",
x"301001000",
x"400301080",
x"520001088",
x"601001000",
x"712002000",
x"801001000",
x"910001008",
x"A01001000",
x"B11002000",
x"C10001001",
x"001001000",
x"046304000",
x"146304000",
x"223302000",
x"301001000",
x"401301020",
x"520001028",
x"601001000",
x"712002000",
x"801001000",
x"910001008",
x"A01001000",
x"B11002000",
x"C10001004",
x"001001000",
x"057504000",
x"157504000",
x"222502000",
x"301001000",
x"400501040",
x"520001048",
x"601001000",
x"724002000",
x"801001000",
x"910001008",
x"A01001000",
x"700001200",
x"B11002000",
x"C10001002",
x"001001000",
x"058404000",
x"158404000",
x"236402000",
x"301001000",
x"400501040",
x"510001048",
x"520001048",
x"601001000",
x"200001100",
x"712002000",
x"801001000",
x"910001008",
x"A01001000",
x"B11002000",
x"C10001002",
x"001001000",
x"057304000",
x"157304000",
x"224302000",
x"301001000",
x"402301010",
x"520001018",
x"601001000",
x"724002000",
x"801001000",
x"910001008",
x"A01001000",
x"700001200",
x"B11002000",
x"C10001001",
x"001001000",
x"045300000",
x"045304000",
x"045304000",
x"045504000",
x"045504000",
x"045504000",
x"046304000",
x"046304000",
x"046304000",
x"047304000",
x"047304000",
x"047304000",
x"145304000",
x"145304000",
x"145304000",
x"145504000",
x"145504000",
x"145504000",
x"146304000",
x"146304000",
x"146304000",
x"147304000",
x"147304000",
x"147304000",
x"222302000",
x"222302000",
x"222302000",
x"222502000",
x"222502000",
x"222502000",
x"223302000",
x"223302000",
x"223302000",
x"224302000",
x"224302000",
x"224302000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"400301080",
x"400301080",
x"400301080",
x"400501040",
x"400501040",
x"400501040",
x"401301020",
x"401301020",
x"401301020",
x"402301010",
x"402301010",
x"402301010",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"C10001004",
x"C10001002",
x"C10001001",
x"C10001004",
x"C10001002",
x"C10001001",
x"C10001004",
x"C10001002",
x"C10001001",
x"C10001004",
x"C10001002",
x"C10001001",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"057304000",
x"057304000",
x"057304000",
x"057504000",
x"057504000",
x"057504000",
x"058304000",
x"058304000",
x"058304000",
x"059304000",
x"059304000",
x"059304000",
x"157304000",
x"157304000",
x"157304000",
x"157504000",
x"157504000",
x"157504000",
x"158304000",
x"158304000",
x"158304000",
x"159304000",
x"159304000",
x"159304000",
x"222302000",
x"222302000",
x"222302000",
x"222502000",
x"222502000",
x"222502000",
x"223302000",
x"223302000",
x"223302000",
x"224302000",
x"224302000",
x"224302000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"400301080",
x"400301080",
x"400301080",
x"400501040",
x"400501040",
x"400501040",
x"401301020",
x"401301020",
x"401301020",
x"402301010",
x"402301010",
x"402301010",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"C10001004",
x"C10001002",
x"C10001001",
x"C10001004",
x"C10001002",
x"C10001001",
x"C10001004",
x"C10001002",
x"C10001001",
x"C10001004",
x"C10001002",
x"C10001001",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"058004000",
x"058004000",
x"058004000",
x"058404000",
x"058404000",
x"058404000",
x"060004000",
x"060004000",
x"060004000",
x"062004000",
x"062004000",
x"062004000",
x"158004000",
x"158004000",
x"158004000",
x"158404000",
x"158404000",
x"158404000",
x"160004000",
x"160004000",
x"160004000",
x"162004000",
x"162004000",
x"162004000",
x"235002000",
x"235002000",
x"235002000",
x"235402000",
x"235402000",
x"235402000",
x"237002000",
x"237002000",
x"237002000",
x"239002000",
x"239002000",
x"239002000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"400301080",
x"400301080",
x"400301080",
x"400501040",
x"400501040",
x"400501040",
x"401301020",
x"401301020",
x"401301020",
x"402301010",
x"402301010",
x"402301010",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"712002000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"C10001008",
x"C10001008",
x"C10001008",
x"C10001008",
x"C10001008",
x"C10001008",
x"C10001008",
x"C10001008",
x"C10001008",
x"C10001008",
x"C10001008",
x"C10001008",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"070004000",
x"070004000",
x"070004000",
x"070404000",
x"070404000",
x"070404000",
x"072004000",
x"072004000",
x"072004000",
x"074004000",
x"074004000",
x"074004000",
x"170004000",
x"170004000",
x"170004000",
x"170404000",
x"170404000",
x"170404000",
x"172004000",
x"172004000",
x"172004000",
x"174004000",
x"174004000",
x"174004000",
x"235002000",
x"235002000",
x"235002000",
x"235002000",
x"235002000",
x"235002000",
x"237002000",
x"237002000",
x"237002000",
x"239002000",
x"239002000",
x"239002000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"301001000",
x"400301080",
x"400301080",
x"400301080",
x"400501040",
x"400501040",
x"400501040",
x"401001020",
x"401001020",
x"401001020",
x"402301010",
x"402301010",
x"402301010",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"510001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"520001008",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"601001000",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"200001100",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"724002000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"801001000",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"910001008",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"A01001000",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"700001200",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"B11002000",
x"C10001004",
x"C10001002",
x"C10001001",
x"C10001004",
x"C10001002",
x"C10001001",
x"C10001004",
x"C10001002",
x"C10001001",
x"C10001004",
x"C10001002",
x"C10001001",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000",
x"001001000"
); 

begin	
process(I)	 
begin 
	case I is
when "0000000000000000000"=> Z <=values(0);  
when "0000100000000100000"=> Z <=values(1);  
when "0000100000000100001"=> Z <=values(2);  
when "0001100000000100001"=> Z <=values(3);  
when "0010100000000100001"=> Z <=values(4);  
when "0011100000000100001"=> Z <=values(5);  
when "0100100000000100001"=> Z <=values(6);  
when "0101100000000100001"=> Z <=values(7);  
when "0110100000000100001"=> Z <=values(8);  
when "0111100000000100001"=> Z <=values(9);  
when "1000100000000100001"=> Z <=values(10); 
when "1001100000000100001"=> Z <=values(11); 
when "1010100000000100001"=> Z <=values(12); 
when "1011100000000100001"=> Z <=values(13); 
when "1100100000000100001"=> Z <=values(14); 
when "0000100000000010000"=> Z <=values(15); 
when "0000100000000010001"=> Z <=values(16); 
when "0001100000000010001"=> Z <=values(17); 
when "0010100000000010001"=> Z <=values(18); 
when "0011100000000010001"=> Z <=values(19); 
when "0100100000000010001"=> Z <=values(20); 
when "0101100000000010001"=> Z <=values(21); 
when "0110100000000010001"=> Z <=values(22); 
when "0111100000000010001"=> Z <=values(23); 
when "1000100000000010001"=> Z <=values(24); 
when "1001100000000010001"=> Z <=values(25); 
when "1010100000000010001"=> Z <=values(26); 
when "1011100000000010001"=> Z <=values(27); 
when "1100100000000010001"=> Z <=values(28); 
when "0000100000000001000"=> Z <=values(29); 
when "0000100000000001001"=> Z <=values(30); 
when "0001100000000001001"=> Z <=values(31); 
when "0010100000000001001"=> Z <=values(32); 
when "0011100000000001001"=> Z <=values(33); 
when "0100100000000001001"=> Z <=values(34); 
when "0101100000000001001"=> Z <=values(35); 
when "0110100000000001001"=> Z <=values(36); 
when "0111100000000001001"=> Z <=values(37); 
when "1000100000000001001"=> Z <=values(38); 
when "1001100000000001001"=> Z <=values(39); 
when "1010100000000001001"=> Z <=values(40); 
when "1010100010000001001"=> Z <=values(41); 
when "1011100000000001001"=> Z <=values(42); 
when "1100100000000001001"=> Z <=values(43); 
when "0000100000000000100"=> Z <=values(44); 
when "0000100000000000101"=> Z <=values(45); 
when "0001100000000000101"=> Z <=values(46); 
when "0010100000000000101"=> Z <=values(47); 
when "0011100000000000101"=> Z <=values(48); 
when "0100100000000000101"=> Z <=values(49); 
when "0100100100000000101"=> Z <=values(50); 
when "0101100000000000101"=> Z <=values(51); 
when "0110100000000000101"=> Z <=values(52); 
when "0110100100000000101"=> Z <=values(53); 
when "0111100000000000101"=> Z <=values(54); 
when "1000100000000000101"=> Z <=values(55); 
when "1001100000000000101"=> Z <=values(56); 
when "1010100000000000101"=> Z <=values(57); 
when "1011100000000000101"=> Z <=values(58); 
when "1100100000000000101"=> Z <=values(59); 
when "0000100000000000010"=> Z <=values(60); 
when "0000100000000000011"=> Z <=values(61); 
when "0001100000000000011"=> Z <=values(62); 
when "0010100000000000011"=> Z <=values(63); 
when "0011100000000000011"=> Z <=values(64); 
when "0100100000000000011"=> Z <=values(65); 
when "0101100000000000011"=> Z <=values(66); 
when "0110100000000000011"=> Z <=values(67); 
when "0111100000000000011"=> Z <=values(68); 
when "1000100000000000011"=> Z <=values(69); 
when "1001100000000000011"=> Z <=values(70); 
when "1010100000000000011"=> Z <=values(71); 
when "1010100010000000011"=> Z <=values(72); 
when "1011100000000000011"=> Z <=values(73); 
when "1100100000000000011"=> Z <=values(74); 
when "0000100000000000000"=> Z <=values(75); 
when "0000100000001000000"=> Z <=values(76); 
when "0000100000010000000"=> Z <=values(77); 
when "0000100000100000000"=> Z <=values(78); 
when "0000100000101000000"=> Z <=values(79); 
when "0000100000110000000"=> Z <=values(80); 
when "0000100001000000000"=> Z <=values(81); 
when "0000100001001000000"=> Z <=values(82); 
when "0000100001010000000"=> Z <=values(83); 
when "0000100001100000000"=> Z <=values(84); 
when "0000100001101000000"=> Z <=values(85); 
when "0000100001110000000"=> Z <=values(86); 
when "0000100000000000001"=> Z <=values(87); 
when "0000100000001000001"=> Z <=values(88); 
when "0000100000010000001"=> Z <=values(89); 
when "0000100000100000001"=> Z <=values(90); 
when "0000100000101000001"=> Z <=values(91); 
when "0000100000110000001"=> Z <=values(92); 
when "0000100001000000001"=> Z <=values(93); 
when "0000100001001000001"=> Z <=values(94); 
when "0000100001010000001"=> Z <=values(95); 
when "0000100001100000001"=> Z <=values(96); 
when "0000100001101000001"=> Z <=values(97); 
when "0000100001110000001"=> Z <=values(98); 
when "0001100000000000001"=> Z <=values(99); 
when "0001100000001000001"=> Z <=values(100);
when "0001100000010000001"=> Z <=values(101);
when "0001100000100000001"=> Z <=values(102);
when "0001100000101000001"=> Z <=values(103);
when "0001100000110000001"=> Z <=values(104);
when "0001100001000000001"=> Z <=values(105);
when "0001100001001000001"=> Z <=values(106);
when "0001100001010000001"=> Z <=values(107);
when "0001100001100000001"=> Z <=values(108);
when "0001100001101000001"=> Z <=values(109);
when "0001100001110000001"=> Z <=values(110);
when "0010100000000000001"=> Z <=values(111);
when "0010100000001000001"=> Z <=values(112);
when "0010100000010000001"=> Z <=values(113);
when "0010100000100000001"=> Z <=values(114);
when "0010100000101000001"=> Z <=values(115);
when "0010100000110000001"=> Z <=values(116);
when "0010100001000000001"=> Z <=values(117);
when "0010100001001000001"=> Z <=values(118);
when "0010100001010000001"=> Z <=values(119);
when "0010100001100000001"=> Z <=values(120);
when "0010100001101000001"=> Z <=values(121);
when "0010100001110000001"=> Z <=values(122);
when "0011100000000000001"=> Z <=values(123);
when "0011100000001000001"=> Z <=values(124);
when "0011100000010000001"=> Z <=values(125);
when "0011100000100000001"=> Z <=values(126);
when "0011100000101000001"=> Z <=values(127);
when "0011100000110000001"=> Z <=values(128);
when "0011100001000000001"=> Z <=values(129);
when "0011100001001000001"=> Z <=values(130);
when "0011100001010000001"=> Z <=values(131);
when "0011100001100000001"=> Z <=values(132);
when "0011100001101000001"=> Z <=values(133);
when "0011100001110000001"=> Z <=values(134);
when "0100100000000000001"=> Z <=values(135);
when "0100100000001000001"=> Z <=values(136);
when "0100100000010000001"=> Z <=values(137);
when "0100100000100000001"=> Z <=values(138);
when "0100100000101000001"=> Z <=values(139);
when "0100100000110000001"=> Z <=values(140);
when "0100100001000000001"=> Z <=values(141);
when "0100100001001000001"=> Z <=values(142);
when "0100100001010000001"=> Z <=values(143);
when "0100100001100000001"=> Z <=values(144);
when "0100100001101000001"=> Z <=values(145);
when "0100100001110000001"=> Z <=values(146);
when "0101100000000000001"=> Z <=values(147);
when "0101100000001000001"=> Z <=values(148);
when "0101100000010000001"=> Z <=values(149);
when "0101100000100000001"=> Z <=values(150);
when "0101100000101000001"=> Z <=values(151);
when "0101100000110000001"=> Z <=values(152);
when "0101100001000000001"=> Z <=values(153);
when "0101100001001000001"=> Z <=values(154);
when "0101100001010000001"=> Z <=values(155);
when "0101100001100000001"=> Z <=values(156);
when "0101100001101000001"=> Z <=values(157);
when "0101100001110000001"=> Z <=values(158);
when "0110100000000000001"=> Z <=values(159);
when "0110100000001000001"=> Z <=values(160);
when "0110100000010000001"=> Z <=values(161);
when "0110100000100000001"=> Z <=values(162);
when "0110100000101000001"=> Z <=values(163);
when "0110100000110000001"=> Z <=values(164);
when "0110100001000000001"=> Z <=values(165);
when "0110100001001000001"=> Z <=values(166);
when "0110100001010000001"=> Z <=values(167);
when "0110100001100000001"=> Z <=values(168);
when "0110100001101000001"=> Z <=values(169);
when "0110100001110000001"=> Z <=values(170);
when "0111100000000000001"=> Z <=values(171);
when "0111100000001000001"=> Z <=values(172);
when "0111100000010000001"=> Z <=values(173);
when "0111100000100000001"=> Z <=values(174);
when "0111100000101000001"=> Z <=values(175);
when "0111100000110000001"=> Z <=values(176);
when "0111100001000000001"=> Z <=values(177);
when "0111100001001000001"=> Z <=values(178);
when "0111100001010000001"=> Z <=values(179);
when "0111100001100000001"=> Z <=values(180);
when "0111100001101000001"=> Z <=values(181);
when "0111100001110000001"=> Z <=values(182);
when "1000100000000000001"=> Z <=values(183);
when "1000100000001000001"=> Z <=values(184);
when "1000100000010000001"=> Z <=values(185);
when "1000100000100000001"=> Z <=values(186);
when "1000100000101000001"=> Z <=values(187);
when "1000100000110000001"=> Z <=values(188);
when "1000100001000000001"=> Z <=values(189);
when "1000100001001000001"=> Z <=values(190);
when "1000100001010000001"=> Z <=values(191);
when "1000100001100000001"=> Z <=values(192);
when "1000100001101000001"=> Z <=values(193);
when "1000100001110000001"=> Z <=values(194);
when "1001100000000000001"=> Z <=values(195);
when "1001100000001000001"=> Z <=values(196);
when "1001100000010000001"=> Z <=values(197);
when "1001100000100000001"=> Z <=values(198);
when "1001100000101000001"=> Z <=values(199);
when "1001100000110000001"=> Z <=values(200);
when "1001100001000000001"=> Z <=values(201);
when "1001100001001000001"=> Z <=values(202);
when "1001100001010000001"=> Z <=values(203);
when "1001100001100000001"=> Z <=values(204);
when "1001100001101000001"=> Z <=values(205);
when "1001100001110000001"=> Z <=values(206);
when "1010100000000000001"=> Z <=values(207);
when "1010100000001000001"=> Z <=values(208);
when "1010100000010000001"=> Z <=values(209);
when "1010100000100000001"=> Z <=values(210);
when "1010100000101000001"=> Z <=values(211);
when "1010100000110000001"=> Z <=values(212);
when "1010100001000000001"=> Z <=values(213);
when "1010100001001000001"=> Z <=values(214);
when "1010100001010000001"=> Z <=values(215);
when "1010100001100000001"=> Z <=values(216);
when "1010100001101000001"=> Z <=values(217);
when "1010100001110000001"=> Z <=values(218);
when "1011100000000000001"=> Z <=values(219);
when "1011100000001000001"=> Z <=values(220);
when "1011100000010000001"=> Z <=values(221);
when "1011100000100000001"=> Z <=values(222);
when "1011100000101000001"=> Z <=values(223);
when "1011100000110000001"=> Z <=values(224);
when "1011100001000000001"=> Z <=values(225);
when "1011100001001000001"=> Z <=values(226);
when "1011100001010000001"=> Z <=values(227);
when "1011100001100000001"=> Z <=values(228);
when "1011100001101000001"=> Z <=values(229);
when "1011100001110000001"=> Z <=values(230);
when "1100100000000000001"=> Z <=values(231);
when "1100100000001000001"=> Z <=values(232);
when "1100100000010000001"=> Z <=values(233);
when "1100100000100000001"=> Z <=values(234);
when "1100100000101000001"=> Z <=values(235);
when "1100100000110000001"=> Z <=values(236);
when "1100100001000000001"=> Z <=values(237);
when "1100100001001000001"=> Z <=values(238);
when "1100100001010000001"=> Z <=values(239);
when "1100100001100000001"=> Z <=values(240);
when "1100100001101000001"=> Z <=values(241);
when "1100100001110000001"=> Z <=values(242);
when "0000101000000000000"=> Z <=values(243);
when "0000101000001000000"=> Z <=values(244);
when "0000101000010000000"=> Z <=values(245);
when "0000101000100000000"=> Z <=values(246);
when "0000101000101000000"=> Z <=values(247);
when "0000101000110000000"=> Z <=values(248);
when "0000101001000000000"=> Z <=values(249);
when "0000101001001000000"=> Z <=values(250);
when "0000101001010000000"=> Z <=values(251);
when "0000101001100000000"=> Z <=values(252);
when "0000101001101000000"=> Z <=values(253);
when "0000101001110000000"=> Z <=values(254);
when "0000101000000000001"=> Z <=values(255);
when "0000101000001000001"=> Z <=values(256);
when "0000101000010000001"=> Z <=values(257);
when "0000101000100000001"=> Z <=values(258);
when "0000101000101000001"=> Z <=values(259);
when "0000101000110000001"=> Z <=values(260);
when "0000101001000000001"=> Z <=values(261);
when "0000101001001000001"=> Z <=values(262);
when "0000101001010000001"=> Z <=values(263);
when "0000101001100000001"=> Z <=values(264);
when "0000101001101000001"=> Z <=values(265);
when "0000101001110000001"=> Z <=values(266);
when "0001101000000000001"=> Z <=values(267);
when "0001101000001000001"=> Z <=values(268);
when "0001101000010000001"=> Z <=values(269);
when "0001101000100000001"=> Z <=values(270);
when "0001101000101000001"=> Z <=values(271);
when "0001101000110000001"=> Z <=values(272);
when "0001101001000000001"=> Z <=values(273);
when "0001101001001000001"=> Z <=values(274);
when "0001101001010000001"=> Z <=values(275);
when "0001101001100000001"=> Z <=values(276);
when "0001101001101000001"=> Z <=values(277);
when "0001101001110000001"=> Z <=values(278);
when "0010101000000000001"=> Z <=values(279);
when "0010101000001000001"=> Z <=values(280);
when "0010101000010000001"=> Z <=values(281);
when "0010101000100000001"=> Z <=values(282);
when "0010101000101000001"=> Z <=values(283);
when "0010101000110000001"=> Z <=values(284);
when "0010101001000000001"=> Z <=values(285);
when "0010101001001000001"=> Z <=values(286);
when "0010101001010000001"=> Z <=values(287);
when "0010101001100000001"=> Z <=values(288);
when "0010101001101000001"=> Z <=values(289);
when "0010101001110000001"=> Z <=values(290);
when "0011101000000000001"=> Z <=values(291);
when "0011101000001000001"=> Z <=values(292);
when "0011101000010000001"=> Z <=values(293);
when "0011101000100000001"=> Z <=values(294);
when "0011101000101000001"=> Z <=values(295);
when "0011101000110000001"=> Z <=values(296);
when "0011101001000000001"=> Z <=values(297);
when "0011101001001000001"=> Z <=values(298);
when "0011101001010000001"=> Z <=values(299);
when "0011101001100000001"=> Z <=values(300);
when "0011101001101000001"=> Z <=values(301);
when "0011101001110000001"=> Z <=values(302);
when "0100101000000000001"=> Z <=values(303);
when "0100101000001000001"=> Z <=values(304);
when "0100101000010000001"=> Z <=values(305);
when "0100101000100000001"=> Z <=values(306);
when "0100101000101000001"=> Z <=values(307);
when "0100101000110000001"=> Z <=values(308);
when "0100101001000000001"=> Z <=values(309);
when "0100101001001000001"=> Z <=values(310);
when "0100101001010000001"=> Z <=values(311);
when "0100101001100000001"=> Z <=values(312);
when "0100101001101000001"=> Z <=values(313);
when "0100101001110000001"=> Z <=values(314);
when "0101101000000000001"=> Z <=values(315);
when "0101101000001000001"=> Z <=values(316);
when "0101101000010000001"=> Z <=values(317);
when "0101101000100000001"=> Z <=values(318);
when "0101101000101000001"=> Z <=values(319);
when "0101101000110000001"=> Z <=values(320);
when "0101101001000000001"=> Z <=values(321);
when "0101101001001000001"=> Z <=values(322);
when "0101101001010000001"=> Z <=values(323);
when "0101101001100000001"=> Z <=values(324);
when "0101101001101000001"=> Z <=values(325);
when "0101101001110000001"=> Z <=values(326);
when "0110101000000000001"=> Z <=values(327);
when "0110101000001000001"=> Z <=values(328);
when "0110101000010000001"=> Z <=values(329);
when "0110101000100000001"=> Z <=values(330);
when "0110101000101000001"=> Z <=values(331);
when "0110101000110000001"=> Z <=values(332);
when "0110101001000000001"=> Z <=values(333);
when "0110101001001000001"=> Z <=values(334);
when "0110101001010000001"=> Z <=values(335);
when "0110101001100000001"=> Z <=values(336);
when "0110101001101000001"=> Z <=values(337);
when "0110101001110000001"=> Z <=values(338);
when "0111101000000000001"=> Z <=values(339);
when "0111101000001000001"=> Z <=values(340);
when "0111101000010000001"=> Z <=values(341);
when "0111101000100000001"=> Z <=values(342);
when "0111101000101000001"=> Z <=values(343);
when "0111101000110000001"=> Z <=values(344);
when "0111101001000000001"=> Z <=values(345);
when "0111101001001000001"=> Z <=values(346);
when "0111101001010000001"=> Z <=values(347);
when "0111101001100000001"=> Z <=values(348);
when "0111101001101000001"=> Z <=values(349);
when "0111101001110000001"=> Z <=values(350);
when "1000101000000000001"=> Z <=values(351);
when "1000101000001000001"=> Z <=values(352);
when "1000101000010000001"=> Z <=values(353);
when "1000101000100000001"=> Z <=values(354);
when "1000101000101000001"=> Z <=values(355);
when "1000101000110000001"=> Z <=values(356);
when "1000101001000000001"=> Z <=values(357);
when "1000101001001000001"=> Z <=values(358);
when "1000101001010000001"=> Z <=values(359);
when "1000101001100000001"=> Z <=values(360);
when "1000101001101000001"=> Z <=values(361);
when "1000101001110000001"=> Z <=values(362);
when "1001101000000000001"=> Z <=values(363);
when "1001101000001000001"=> Z <=values(364);
when "1001101000010000001"=> Z <=values(365);
when "1001101000100000001"=> Z <=values(366);
when "1001101000101000001"=> Z <=values(367);
when "1001101000110000001"=> Z <=values(368);
when "1001101001000000001"=> Z <=values(369);
when "1001101001001000001"=> Z <=values(370);
when "1001101001010000001"=> Z <=values(371);
when "1001101001100000001"=> Z <=values(372);
when "1001101001101000001"=> Z <=values(373);
when "1001101001110000001"=> Z <=values(374);
when "1010101000000000001"=> Z <=values(375);
when "1010101000001000001"=> Z <=values(376);
when "1010101000010000001"=> Z <=values(377);
when "1010101000100000001"=> Z <=values(378);
when "1010101000101000001"=> Z <=values(379);
when "1010101000110000001"=> Z <=values(380);
when "1010101001000000001"=> Z <=values(381);
when "1010101001001000001"=> Z <=values(382);
when "1010101001010000001"=> Z <=values(383);
when "1010101001100000001"=> Z <=values(384);
when "1010101001101000001"=> Z <=values(385);
when "1010101001110000001"=> Z <=values(386);
when "1010101010000000001"=> Z <=values(387);
when "1010101010001000001"=> Z <=values(388);
when "1010101010010000001"=> Z <=values(389);
when "1010101010100000001"=> Z <=values(390);
when "1010101010101000001"=> Z <=values(391);
when "1010101010110000001"=> Z <=values(392);
when "1010101011000000001"=> Z <=values(393);
when "1010101011001000001"=> Z <=values(394);
when "1010101011010000001"=> Z <=values(395);
when "1010101011100000001"=> Z <=values(396);
when "1010101011101000001"=> Z <=values(397);
when "1010101011110000001"=> Z <=values(398);
when "1011101000000000001"=> Z <=values(399);
when "1011101000001000001"=> Z <=values(400);
when "1011101000010000001"=> Z <=values(401);
when "1011101000100000001"=> Z <=values(402);
when "1011101000101000001"=> Z <=values(403);
when "1011101000110000001"=> Z <=values(404);
when "1011101001000000001"=> Z <=values(405);
when "1011101001001000001"=> Z <=values(406);
when "1011101001010000001"=> Z <=values(407);
when "1011101001100000001"=> Z <=values(408);
when "1011101001101000001"=> Z <=values(409);
when "1011101001110000001"=> Z <=values(410);
when "1100101000000000001"=> Z <=values(411);
when "1100101000001000001"=> Z <=values(412);
when "1100101000010000001"=> Z <=values(413);
when "1100101000100000001"=> Z <=values(414);
when "1100101000101000001"=> Z <=values(415);
when "1100101000110000001"=> Z <=values(416);
when "1100101001000000001"=> Z <=values(417);
when "1100101001001000001"=> Z <=values(418);
when "1100101001010000001"=> Z <=values(419);
when "1100101001100000001"=> Z <=values(420);
when "1100101001101000001"=> Z <=values(421);
when "1100101001110000001"=> Z <=values(422);
when "0000110000000000000"=> Z <=values(423);
when "0000110000001000000"=> Z <=values(424);
when "0000110000010000000"=> Z <=values(425);
when "0000110000100000000"=> Z <=values(426);
when "0000110000101000000"=> Z <=values(427);
when "0000110000110000000"=> Z <=values(428);
when "0000110001000000000"=> Z <=values(429);
when "0000110001001000000"=> Z <=values(430);
when "0000110001010000000"=> Z <=values(431);
when "0000110001100000000"=> Z <=values(432);
when "0000110001101000000"=> Z <=values(433);
when "0000110001110000000"=> Z <=values(434);
when "0000110000000000001"=> Z <=values(435);
when "0000110000001000001"=> Z <=values(436);
when "0000110000010000001"=> Z <=values(437);
when "0000110000100000001"=> Z <=values(438);
when "0000110000101000001"=> Z <=values(439);
when "0000110000110000001"=> Z <=values(440);
when "0000110001000000001"=> Z <=values(441);
when "0000110001001000001"=> Z <=values(442);
when "0000110001010000001"=> Z <=values(443);
when "0000110001100000001"=> Z <=values(444);
when "0000110001101000001"=> Z <=values(445);
when "0000110001110000001"=> Z <=values(446);
when "0001110000000000001"=> Z <=values(447);
when "0001110000001000001"=> Z <=values(448);
when "0001110000010000001"=> Z <=values(449);
when "0001110000100000001"=> Z <=values(450);
when "0001110000101000001"=> Z <=values(451);
when "0001110000110000001"=> Z <=values(452);
when "0001110001000000001"=> Z <=values(453);
when "0001110001001000001"=> Z <=values(454);
when "0001110001010000001"=> Z <=values(455);
when "0001110001100000001"=> Z <=values(456);
when "0001110001101000001"=> Z <=values(457);
when "0001110001110000001"=> Z <=values(458);
when "0010110000000000001"=> Z <=values(459);
when "0010110000001000001"=> Z <=values(460);
when "0010110000010000001"=> Z <=values(461);
when "0010110000100000001"=> Z <=values(462);
when "0010110000101000001"=> Z <=values(463);
when "0010110000110000001"=> Z <=values(464);
when "0010110001000000001"=> Z <=values(465);
when "0010110001001000001"=> Z <=values(466);
when "0010110001010000001"=> Z <=values(467);
when "0010110001100000001"=> Z <=values(468);
when "0010110001101000001"=> Z <=values(469);
when "0010110001110000001"=> Z <=values(470);
when "0011110000000000001"=> Z <=values(471);
when "0011110000001000001"=> Z <=values(472);
when "0011110000010000001"=> Z <=values(473);
when "0011110000100000001"=> Z <=values(474);
when "0011110000101000001"=> Z <=values(475);
when "0011110000110000001"=> Z <=values(476);
when "0011110001000000001"=> Z <=values(477);
when "0011110001001000001"=> Z <=values(478);
when "0011110001010000001"=> Z <=values(479);
when "0011110001100000001"=> Z <=values(480);
when "0011110001101000001"=> Z <=values(481);
when "0011110001110000001"=> Z <=values(482);
when "0100110000000000001"=> Z <=values(483);
when "0100110000001000001"=> Z <=values(484);
when "0100110000010000001"=> Z <=values(485);
when "0100110000100000001"=> Z <=values(486);
when "0100110000101000001"=> Z <=values(487);
when "0100110000110000001"=> Z <=values(488);
when "0100110001000000001"=> Z <=values(489);
when "0100110001001000001"=> Z <=values(490);
when "0100110001010000001"=> Z <=values(491);
when "0100110001100000001"=> Z <=values(492);
when "0100110001101000001"=> Z <=values(493);
when "0100110001110000001"=> Z <=values(494);
when "0100110100000000001"=> Z <=values(495);
when "0100110100001000001"=> Z <=values(496);
when "0100110100010000001"=> Z <=values(497);
when "0100110100100000001"=> Z <=values(498);
when "0100110100101000001"=> Z <=values(499);
when "0100110100110000001"=> Z <=values(500);
when "0100110101000000001"=> Z <=values(501);
when "0100110101001000001"=> Z <=values(502);
when "0100110101010000001"=> Z <=values(503);
when "0100110101100000001"=> Z <=values(504);
when "0100110101101000001"=> Z <=values(505);
when "0100110101110000001"=> Z <=values(506);
when "0101110000000000001"=> Z <=values(507);
when "0101110000001000001"=> Z <=values(508);
when "0101110000010000001"=> Z <=values(509);
when "0101110000100000001"=> Z <=values(510);
when "0101110000101000001"=> Z <=values(511);
when "0101110000110000001"=> Z <=values(512);
when "0101110001000000001"=> Z <=values(513);
when "0101110001001000001"=> Z <=values(514);
when "0101110001010000001"=> Z <=values(515);
when "0101110001100000001"=> Z <=values(516);
when "0101110001101000001"=> Z <=values(517);
when "0101110001110000001"=> Z <=values(518);
when "0110110000000000001"=> Z <=values(519);
when "0110110000001000001"=> Z <=values(520);
when "0110110000010000001"=> Z <=values(521);
when "0110110000100000001"=> Z <=values(522);
when "0110110000101000001"=> Z <=values(523);
when "0110110000110000001"=> Z <=values(524);
when "0110110001000000001"=> Z <=values(525);
when "0110110001001000001"=> Z <=values(526);
when "0110110001010000001"=> Z <=values(527);
when "0110110001100000001"=> Z <=values(528);
when "0110110001101000001"=> Z <=values(529);
when "0110110001110000001"=> Z <=values(530);
when "0110110100000000001"=> Z <=values(531);
when "0110110100001000001"=> Z <=values(532);
when "0110110100010000001"=> Z <=values(533);
when "0110110100100000001"=> Z <=values(534);
when "0110110100101000001"=> Z <=values(535);
when "0110110100110000001"=> Z <=values(536);
when "0110110101000000001"=> Z <=values(537);
when "0110110101001000001"=> Z <=values(538);
when "0110110101010000001"=> Z <=values(539);
when "0110110101100000001"=> Z <=values(540);
when "0110110101101000001"=> Z <=values(541);
when "0110110101110000001"=> Z <=values(542);
when "0111110000000000001"=> Z <=values(543);
when "0111110000001000001"=> Z <=values(544);
when "0111110000010000001"=> Z <=values(545);
when "0111110000100000001"=> Z <=values(546);
when "0111110000101000001"=> Z <=values(547);
when "0111110000110000001"=> Z <=values(548);
when "0111110001000000001"=> Z <=values(549);
when "0111110001001000001"=> Z <=values(550);
when "0111110001010000001"=> Z <=values(551);
when "0111110001100000001"=> Z <=values(552);
when "0111110001101000001"=> Z <=values(553);
when "0111110001110000001"=> Z <=values(554);
when "1000110000000000001"=> Z <=values(555);
when "1000110000001000001"=> Z <=values(556);
when "1000110000010000001"=> Z <=values(557);
when "1000110000100000001"=> Z <=values(558);
when "1000110000101000001"=> Z <=values(559);
when "1000110000110000001"=> Z <=values(560);
when "1000110001000000001"=> Z <=values(561);
when "1000110001001000001"=> Z <=values(562);
when "1000110001010000001"=> Z <=values(563);
when "1000110001100000001"=> Z <=values(564);
when "1000110001101000001"=> Z <=values(565);
when "1000110001110000001"=> Z <=values(566);
when "1001110000000000001"=> Z <=values(567);
when "1001110000001000001"=> Z <=values(568);
when "1001110000010000001"=> Z <=values(569);
when "1001110000100000001"=> Z <=values(570);
when "1001110000101000001"=> Z <=values(571);
when "1001110000110000001"=> Z <=values(572);
when "1001110001000000001"=> Z <=values(573);
when "1001110001001000001"=> Z <=values(574);
when "1001110001010000001"=> Z <=values(575);
when "1001110001100000001"=> Z <=values(576);
when "1001110001101000001"=> Z <=values(577);
when "1001110001110000001"=> Z <=values(578);
when "1010110000000000001"=> Z <=values(579);
when "1010110000001000001"=> Z <=values(580);
when "1010110000010000001"=> Z <=values(581);
when "1010110000100000001"=> Z <=values(582);
when "1010110000101000001"=> Z <=values(583);
when "1010110000110000001"=> Z <=values(584);
when "1010110001000000001"=> Z <=values(585);
when "1010110001001000001"=> Z <=values(586);
when "1010110001010000001"=> Z <=values(587);
when "1010110001100000001"=> Z <=values(588);
when "1010110001101000001"=> Z <=values(589);
when "1010110001110000001"=> Z <=values(590);
when "1011110000000000001"=> Z <=values(591);
when "1011110000001000001"=> Z <=values(592);
when "1011110000010000001"=> Z <=values(593);
when "1011110000100000001"=> Z <=values(594);
when "1011110000101000001"=> Z <=values(595);
when "1011110000110000001"=> Z <=values(596);
when "1011110001000000001"=> Z <=values(597);
when "1011110001001000001"=> Z <=values(598);
when "1011110001010000001"=> Z <=values(599);
when "1011110001100000001"=> Z <=values(600);
when "1011110001101000001"=> Z <=values(601);
when "1011110001110000001"=> Z <=values(602);
when "1100110000000000001"=> Z <=values(603);
when "1100110000001000001"=> Z <=values(604);
when "1100110000010000001"=> Z <=values(605);
when "1100110000100000001"=> Z <=values(606);
when "1100110000101000001"=> Z <=values(607);
when "1100110000110000001"=> Z <=values(608);
when "1100110001000000001"=> Z <=values(609);
when "1100110001001000001"=> Z <=values(610);
when "1100110001010000001"=> Z <=values(611);
when "1100110001100000001"=> Z <=values(612);
when "1100110001101000001"=> Z <=values(613);
when "1100110001110000001"=> Z <=values(614);
when "0000111000000000000"=> Z <=values(615);
when "0000111000001000000"=> Z <=values(616);
when "0000111000010000000"=> Z <=values(617);
when "0000111000100000000"=> Z <=values(618);
when "0000111000101000000"=> Z <=values(619);
when "0000111000110000000"=> Z <=values(620);
when "0000111001000000000"=> Z <=values(621);
when "0000111001001000000"=> Z <=values(622);
when "0000111001010000000"=> Z <=values(623);
when "0000111001100000000"=> Z <=values(624);
when "0000111001101000000"=> Z <=values(625);
when "0000111001110000000"=> Z <=values(626);
when "0000111000000000001"=> Z <=values(627);
when "0000111000001000001"=> Z <=values(628);
when "0000111000010000001"=> Z <=values(629);
when "0000111000100000001"=> Z <=values(630);
when "0000111000101000001"=> Z <=values(631);
when "0000111000110000001"=> Z <=values(632);
when "0000111001000000001"=> Z <=values(633);
when "0000111001001000001"=> Z <=values(634);
when "0000111001010000001"=> Z <=values(635);
when "0000111001100000001"=> Z <=values(636);
when "0000111001101000001"=> Z <=values(637);
when "0000111001110000001"=> Z <=values(638);
when "0001111000000000001"=> Z <=values(639);
when "0001111000001000001"=> Z <=values(640);
when "0001111000010000001"=> Z <=values(641);
when "0001111000100000001"=> Z <=values(642);
when "0001111000101000001"=> Z <=values(643);
when "0001111000110000001"=> Z <=values(644);
when "0001111001000000001"=> Z <=values(645);
when "0001111001001000001"=> Z <=values(646);
when "0001111001010000001"=> Z <=values(647);
when "0001111001100000001"=> Z <=values(648);
when "0001111001101000001"=> Z <=values(649);
when "0001111001110000001"=> Z <=values(650);
when "0010111000000000001"=> Z <=values(651);
when "0010111000001000001"=> Z <=values(652);
when "0010111000010000001"=> Z <=values(653);
when "0010111000100000001"=> Z <=values(654);
when "0010111000101000001"=> Z <=values(655);
when "0010111000110000001"=> Z <=values(656);
when "0010111001000000001"=> Z <=values(657);
when "0010111001001000001"=> Z <=values(658);
when "0010111001010000001"=> Z <=values(659);
when "0010111001100000001"=> Z <=values(660);
when "0010111001101000001"=> Z <=values(661);
when "0010111001110000001"=> Z <=values(662);
when "0011111000000000001"=> Z <=values(663);
when "0011111000001000001"=> Z <=values(664);
when "0011111000010000001"=> Z <=values(665);
when "0011111000100000001"=> Z <=values(666);
when "0011111000101000001"=> Z <=values(667);
when "0011111000110000001"=> Z <=values(668);
when "0011111001000000001"=> Z <=values(669);
when "0011111001001000001"=> Z <=values(670);
when "0011111001010000001"=> Z <=values(671);
when "0011111001100000001"=> Z <=values(672);
when "0011111001101000001"=> Z <=values(673);
when "0011111001110000001"=> Z <=values(674);
when "0100111000000000001"=> Z <=values(675);
when "0100111000001000001"=> Z <=values(676);
when "0100111000010000001"=> Z <=values(677);
when "0100111000100000001"=> Z <=values(678);
when "0100111000101000001"=> Z <=values(679);
when "0100111000110000001"=> Z <=values(680);
when "0100111001000000001"=> Z <=values(681);
when "0100111001001000001"=> Z <=values(682);
when "0100111001010000001"=> Z <=values(683);
when "0100111001100000001"=> Z <=values(684);
when "0100111001101000001"=> Z <=values(685);
when "0100111001110000001"=> Z <=values(686);
when "0100111100000000001"=> Z <=values(687);
when "0100111100001000001"=> Z <=values(688);
when "0100111100010000001"=> Z <=values(689);
when "0100111100100000001"=> Z <=values(690);
when "0100111100101000001"=> Z <=values(691);
when "0100111100110000001"=> Z <=values(692);
when "0100111101000000001"=> Z <=values(693);
when "0100111101001000001"=> Z <=values(694);
when "0100111101010000001"=> Z <=values(695);
when "0100111101100000001"=> Z <=values(696);
when "0100111101101000001"=> Z <=values(697);
when "0100111101110000001"=> Z <=values(698);
when "0101111000000000001"=> Z <=values(699);
when "0101111000001000001"=> Z <=values(700);
when "0101111000010000001"=> Z <=values(701);
when "0101111000100000001"=> Z <=values(702);
when "0101111000101000001"=> Z <=values(703);
when "0101111000110000001"=> Z <=values(704);
when "0101111001000000001"=> Z <=values(705);
when "0101111001001000001"=> Z <=values(706);
when "0101111001010000001"=> Z <=values(707);
when "0101111001100000001"=> Z <=values(708);
when "0101111001101000001"=> Z <=values(709);
when "0101111001110000001"=> Z <=values(710);
when "0110111000000000001"=> Z <=values(711);
when "0110111000001000001"=> Z <=values(712);
when "0110111000010000001"=> Z <=values(713);
when "0110111000100000001"=> Z <=values(714);
when "0110111000101000001"=> Z <=values(715);
when "0110111000110000001"=> Z <=values(716);
when "0110111001000000001"=> Z <=values(717);
when "0110111001001000001"=> Z <=values(718);
when "0110111001010000001"=> Z <=values(719);
when "0110111001100000001"=> Z <=values(720);
when "0110111001101000001"=> Z <=values(721);
when "0110111001110000001"=> Z <=values(722);
when "0110111100000000001"=> Z <=values(723);
when "0110111100001000001"=> Z <=values(724);
when "0110111100010000001"=> Z <=values(725);
when "0110111100100000001"=> Z <=values(726);
when "0110111100101000001"=> Z <=values(727);
when "0110111100110000001"=> Z <=values(728);
when "0110111101000000001"=> Z <=values(729);
when "0110111101001000001"=> Z <=values(730);
when "0110111101010000001"=> Z <=values(731);
when "0110111101100000001"=> Z <=values(732);
when "0110111101101000001"=> Z <=values(733);
when "0110111101110000001"=> Z <=values(734);
when "0111111000000000001"=> Z <=values(735);
when "0111111000001000001"=> Z <=values(736);
when "0111111000010000001"=> Z <=values(737);
when "0111111000100000001"=> Z <=values(738);
when "0111111000101000001"=> Z <=values(739);
when "0111111000110000001"=> Z <=values(740);
when "0111111001000000001"=> Z <=values(741);
when "0111111001001000001"=> Z <=values(742);
when "0111111001010000001"=> Z <=values(743);
when "0111111001100000001"=> Z <=values(744);
when "0111111001101000001"=> Z <=values(745);
when "0111111001110000001"=> Z <=values(746);
when "1000111000000000001"=> Z <=values(747);
when "1000111000001000001"=> Z <=values(748);
when "1000111000010000001"=> Z <=values(749);
when "1000111000100000001"=> Z <=values(750);
when "1000111000101000001"=> Z <=values(751);
when "1000111000110000001"=> Z <=values(752);
when "1000111001000000001"=> Z <=values(753);
when "1000111001001000001"=> Z <=values(754);
when "1000111001010000001"=> Z <=values(755);
when "1000111001100000001"=> Z <=values(756);
when "1000111001101000001"=> Z <=values(757);
when "1000111001110000001"=> Z <=values(758);
when "1001111000000000001"=> Z <=values(759);
when "1001111000001000001"=> Z <=values(760);
when "1001111000010000001"=> Z <=values(761);
when "1001111000100000001"=> Z <=values(762);
when "1001111000101000001"=> Z <=values(763);
when "1001111000110000001"=> Z <=values(764);
when "1001111001000000001"=> Z <=values(765);
when "1001111001001000001"=> Z <=values(766);
when "1001111001010000001"=> Z <=values(767);
when "1001111001100000001"=> Z <=values(768);
when "1001111001101000001"=> Z <=values(769);
when "1001111001110000001"=> Z <=values(770);
when "1010111000000000001"=> Z <=values(771);
when "1010111000001000001"=> Z <=values(772);
when "1010111000010000001"=> Z <=values(773);
when "1010111000100000001"=> Z <=values(774);
when "1010111000101000001"=> Z <=values(775);
when "1010111000110000001"=> Z <=values(776);
when "1010111001000000001"=> Z <=values(777);
when "1010111001001000001"=> Z <=values(778);
when "1010111001010000001"=> Z <=values(779);
when "1010111001100000001"=> Z <=values(780);
when "1010111001101000001"=> Z <=values(781);
when "1010111001110000001"=> Z <=values(782);
when "1010111010000000001"=> Z <=values(783);
when "1010111010001000001"=> Z <=values(784);
when "1010111010010000001"=> Z <=values(785);
when "1010111010100000001"=> Z <=values(786);
when "1010111010101000001"=> Z <=values(787);
when "1010111010110000001"=> Z <=values(788);
when "1010111011000000001"=> Z <=values(789);
when "1010111011001000001"=> Z <=values(790);
when "1010111011010000001"=> Z <=values(791);
when "1010111011100000001"=> Z <=values(792);
when "1010111011101000001"=> Z <=values(793);
when "1010111011110000001"=> Z <=values(794);
when "1011111000000000001"=> Z <=values(795);
when "1011111000001000001"=> Z <=values(796);
when "1011111000010000001"=> Z <=values(797);
when "1011111000100000001"=> Z <=values(798);
when "1011111000101000001"=> Z <=values(799);
when "1011111000110000001"=> Z <=values(800);
when "1011111001000000001"=> Z <=values(801);
when "1011111001001000001"=> Z <=values(802);
when "1011111001010000001"=> Z <=values(803);
when "1011111001100000001"=> Z <=values(804);
when "1011111001101000001"=> Z <=values(805);
when "1011111001110000001"=> Z <=values(806);
when "1100111000000000001"=> Z <=values(807);
when "1100111000001000001"=> Z <=values(808);
when "1100111000010000001"=> Z <=values(809);
when "1100111000100000001"=> Z <=values(810);
when "1100111000101000001"=> Z <=values(811);
when "1100111000110000001"=> Z <=values(812);
when "1100111001000000001"=> Z <=values(813);
when "1100111001001000001"=> Z <=values(814);
when "1100111001010000001"=> Z <=values(815);
when "1100111001100000001"=> Z <=values(816);
when "1100111001101000001"=> Z <=values(817);
when "1100111001110000001"=> Z <=values(818);	
		when others => Z <=(x"000000000");
	end case; 
end process;

	

end ROM_WASH;
